*IV CHARACTERISTICS
Vgs vgs 0 0
Vds vds 0 -1.8

M1 vds vgs 0 0 PMOS L=60n W={W}
.model PMOS PMOS
.dc Vgs 0 -5 -0.1
.step param W 120n 480n 120n
.backanno
.end
